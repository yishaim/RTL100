`timescale 1ns / 1ps

//Day 1 - 2 to 1 mux with 8 bit inputs and output

module top(
    input wire [7:0] a_i,
    input wire [7:0] b_i,
    input wire sel_i,
    output wire [7:0] y_o
    );
    
    assign y_o = sel_i ? a_i : b_i;
    
   
endmodule
